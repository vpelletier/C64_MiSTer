// 
// c1541_track
// Copyright (c) 2016 Sorgelig
//
// This source file is free software: you can redistribute it and/or modify
// it under the terms of the Lesser GNU General Public License as published
// by the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
//
// This source file is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <http://www.gnu.org/licenses/>.
//
//
/////////////////////////////////////////////////////////////////////////

module c1541_track
(
	input         clk,
	input         reset,

	input         sd_clk,
	output [31:0] sd_lba,
	output reg    sd_rd,
	output reg    sd_wr,
	input         sd_ack,

	input   [8:0] sd_buff_addr,
	input   [7:0] sd_buff_dout,
	output  [7:0] sd_buff_din,
	input         sd_buff_wr,

	input         disk_change,
	input   [1:0] stp,
	input         mtr,
	input         act,
	output reg    tr00_sense_n,
	output reg    buff_dout,
	input         buff_din,
	input         buff_we,
	output reg    busy
);

always @(posedge sd_clk) begin
	reg wr1,rd1;
	
	wr1 <= wr;
	rd1 <= rd;
	
	sd_wr <= wr1;
	sd_rd <= rd1;
end

wire [62:0] rnd;
lfsr random(rnd);

assign sd_buff_din = ~metadata_track ? sd_track_buff_din :
		     sd_buff_addr[1:0] == 2'b00 ? sd_metadata_buff_din[31:24] :
		     sd_buff_addr[1:0] == 2'b01 ? sd_metadata_buff_din[23:16] :
		     sd_buff_addr[1:0] == 2'b10 ? sd_metadata_buff_din[15: 8] :
						  sd_metadata_buff_din[ 7: 0];

wire sd_b_ack = sd_ack & busy;
reg [15:0] buff_bit_addr;
wire [15:0] next_buff_bit_addr = buff_bit_addr + 16'b1;
wire [7:0] buff_dout_byte;
wire flux_change = buff_dout_byte[~buff_bit_addr[2:0]];
wire buff_din_posedge = !old_buff_din && buff_din;
reg old_buff_din;
reg buff_din_latched;

wire [7:0] sd_track_buff_din;
wire [7:0] buff_din_byte = buff_bit_addr[2:0] == 3'd0 ? {                     buff_din_latched, buff_dout_byte[6:0]} :
			   buff_bit_addr[2:0] == 3'd1 ? {buff_dout_byte[7  ], buff_din_latched, buff_dout_byte[5:0]} :
			   buff_bit_addr[2:0] == 3'd2 ? {buff_dout_byte[7:6], buff_din_latched, buff_dout_byte[4:0]} :
			   buff_bit_addr[2:0] == 3'd3 ? {buff_dout_byte[7:5], buff_din_latched, buff_dout_byte[3:0]} :
			   buff_bit_addr[2:0] == 3'd4 ? {buff_dout_byte[7:4], buff_din_latched, buff_dout_byte[2:0]} :
			   buff_bit_addr[2:0] == 3'd5 ? {buff_dout_byte[7:3], buff_din_latched, buff_dout_byte[1:0]} :
			   buff_bit_addr[2:0] == 3'd6 ? {buff_dout_byte[7:2], buff_din_latched, buff_dout_byte[  0]} :
							{buff_dout_byte[7:1], buff_din_latched                     };
trk_dpram buffer
(
	.clock_a(sd_clk),
	.address_a({sd_buff_base, sd_buff_addr}),
	.data_a(sd_buff_dout),
	.wren_a(sd_b_ack & sd_buff_wr & ~metadata_track),
	.q_a(sd_track_buff_din),

	.clock_b(clk),
	.address_b(buff_bit_addr[15:3]),
	.data_b(buff_din_byte),
	.wren_b(buff_we),
	.q_b(buff_dout_byte)
);

wire [31:0] sd_metadata_buff_din;
wire [31:0] sd_metadata_buff_dout = sd_buff_addr[1:0] == 2'b00 ? {                             sd_buff_dout, sd_metadata_buff_din[23:0]} :
				    sd_buff_addr[1:0] == 2'b01 ? {sd_metadata_buff_din[31:24], sd_buff_dout, sd_metadata_buff_din[15:0]} :
				    sd_buff_addr[1:0] == 2'b10 ? {sd_metadata_buff_din[31:16], sd_buff_dout, sd_metadata_buff_din[ 7:0]} :
								 {sd_metadata_buff_din[31: 8], sd_buff_dout                            };
wire [1:0] speed_zone;
wire [5:0] delay_integer;
wire [7:0] delay_fractional;
wire [15:0] track_length;

trk_dpram #(.DATAWIDTH(32), .ADDRWIDTH(7)) metadata_buffer
(
	.clock_a(sd_clk),
	.address_a(sd_buff_addr[8:2]),
	.data_a(sd_metadata_buff_dout),
	.wren_a(sd_b_ack & sd_buff_wr & metadata_track),
	.q_a(sd_metadata_buff_din),

	.clock_b(clk),
	.address_b(cur_half_track),
	.data_b(), // XXX: no write support
	.wren_b(1'b0),
	.q_b({speed_zone, delay_integer, delay_fractional, track_length})
);

reg [3:0] sd_buff_base;
reg [6:0] cur_half_track;
wire metadata_track = cur_half_track == 7'd84;
assign sd_lba = {cur_half_track, sd_buff_base};
reg rd,wr;

always @(posedge clk) begin
	reg ack1,ack2,ack;
	reg old_ack;
	reg old_disk_change, ready = 0;
	reg saving = 0;
	reg [62:0] rnd_reg;
	reg [7:0] clk_counter;
	reg [7:0] clk_counter_max_integer;
	reg [7:0] clk_counter_max_fractional;
	reg [1:0] no_flux_change_count;

	old_disk_change <= disk_change;
	if (~old_disk_change && disk_change) ready <= 1;

	old_buff_din <= buff_din;
	if (mtr) begin
		if (clk_counter == clk_counter_max_integer) begin
			{clk_counter_max_integer, clk_counter_max_fractional} <= {1'b0, delay_integer, delay_fractional, 1'b0} + {1'b0, 6'd32, clk_counter_max_fractional, 1'b0};
			buff_bit_addr <= next_buff_bit_addr[15:3] < track_length ? next_buff_bit_addr : 16'b0;
			buff_din_latched <= buff_din_posedge;
			rnd_reg <= rnd;
			clk_counter <= 0;
		end else begin
			if (clk_counter == 6'd1) begin
				if (flux_change) begin
					buff_dout <= ~buff_we;
					no_flux_change_count <= 0;
				end else begin
					// a zero lasts twice as long as a one
					//clk_counter_max_integer <= {clk_counter_max_integer[6:0], 1'b0};
					if (no_flux_change_count == 2'b11) begin
						buff_dout <= ~buff_we & rnd_reg[0];
					end else begin
						buff_dout <= 0;
						no_flux_change_count <= no_flux_change_count + 2'b1;
					end
				end
			end else if (clk_counter == 6'd8)
				buff_dout <= 0;
			buff_din_latched <= buff_din_latched | buff_din_posedge;
			clk_counter <= clk_counter + 6'b1;
		end
	end

	ack1 <= sd_b_ack;
	ack2 <= ack1;
	if(ack2 == ack1) ack <= ack1;

	old_ack <= ack;
	if(ack) {rd,wr} <= 0;

	if(reset) begin
		cur_half_track <= 0;
		busy  <= 0;
		rd <= 0;
		wr <= 0;
		saving<= 0;
	end
	else
	if(busy) begin
		if(old_ack && ~ack) begin
			if(metadata_track) begin
				cur_half_track <= half_track;
				rd <= 1;
			end
			else
			if(sd_buff_base != 4'b1111) begin
				sd_buff_base <= sd_buff_base + 4'b1;
				if(saving) wr <= 1;
					else rd <= 1;
			end
			else
			if(saving && (cur_half_track != half_track)) begin
				saving <= 0;
				cur_half_track <= half_track;
				sd_buff_base <= 0;
				rd <= 1;
			end
			else
			begin
				busy <= 0;
			end
		end
	end
	else
	if(ready) begin
		if(save_track) begin
			saving <= 1;
			sd_buff_base <= 0;
			wr <= 1;
			busy <= 1;
		end
		else
		if (
			(cur_half_track != half_track) ||
			(old_disk_change && ~disk_change)
		) begin
			saving <= 0;
			cur_half_track <= old_disk_change && ~disk_change ? 7'd84 : half_track;
			sd_buff_base <= 0;
			rd <= 1;
			busy <= 1;
		end
	end
end

reg [6:0] half_track;
reg       save_track;
always @(posedge clk) begin
	reg       track_modified;
	reg [1:0] stp_r;
	reg       act_r;

	tr00_sense_n <= |half_track;
	stp_r <= stp;
	act_r <= act;
	save_track <= 0;

	if (buff_we) track_modified <= 1;
	if (disk_change) track_modified <= 0;

	if (reset) begin
		half_track <= 36;
		track_modified <= 0;
	end else begin
		if (mtr) begin
			if ((stp_r == 0 && stp == 1)
				|| (stp_r == 1 && stp == 2)
				|| (stp_r == 2 && stp == 3)
				|| (stp_r == 3 && stp == 0)) begin
				if (half_track < 83) half_track <= half_track + 7'b1;
				save_track <= track_modified;
				track_modified <= 0;
			end

			if ((stp_r == 0 && stp == 3)
				|| (stp_r == 3 && stp == 2)
				|| (stp_r == 2 && stp == 1)
				|| (stp_r == 1 && stp == 0)) begin
				if (half_track) half_track <= half_track - 7'b1;
				save_track <= track_modified;
				track_modified <= 0;
			end
		end

		if (act_r && ~act) begin		// stopping activity
			save_track <= track_modified;
			track_modified <= 0;
		end
	end
end
endmodule

module trk_dpram #(parameter DATAWIDTH=8, ADDRWIDTH=13)
(
	input	                     clock_a,
	input	     [ADDRWIDTH-1:0] address_a,
	input	     [DATAWIDTH-1:0] data_a,
	input	                     wren_a,
	output reg [DATAWIDTH-1:0] q_a,

	input	                     clock_b,
	input	     [ADDRWIDTH-1:0] address_b,
	input	     [DATAWIDTH-1:0] data_b,
	input	                     wren_b,
	output reg [DATAWIDTH-1:0] q_b
);

logic [DATAWIDTH-1:0] ram[0:(1<<ADDRWIDTH)-1];

always_ff@(posedge clock_a) begin
	if(wren_a) begin
		ram[address_a] <= data_a;
		q_a <= data_a;
	end else begin
		q_a <= ram[address_a];
	end
end

always_ff@(posedge clock_b) begin
	if(wren_b) begin
		ram[address_b] <= data_b;
		q_b <= data_b;
	end else begin
		q_b <= ram[address_b];
	end
end

endmodule
